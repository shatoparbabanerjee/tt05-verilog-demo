`default_nettype none

module current_based_tt_um_lif (
    input  wire [7:0] ui_in,    // Dedicated inputs - connected to the input switches
    output wire [7:0] uo_out,   // Dedicated outputs - connected to the 7 segment display
    input  wire [7:0] uio_in,   // IOs: Bidirectional Input path
    output wire [7:0] uio_out,  // IOs: Bidirectional Output path
    output wire [7:0] uio_oe,   // IOs: Bidirectional Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // will go high when the design is enabled
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

    assign uio_oe = 8'b11111111;
    assign uio_out[6:0] = 7'd0;

    wire spike;
    wire [7:0] membrane_potential;

    // Instantiate the current-based LIF neuron
    current_based_lif lif1(.synaptic_current(ui_in), .clk(clk), .rst_n(rst_n), .spike(spike), .membrane_potential(membrane_potential));

    // Connect the LIF neuron output to the 7-segment display output
    assign uo_out = {spike, membrane_potential[6:0]};

endmodule
